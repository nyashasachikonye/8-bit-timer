LIBRARY altera;
USE altera.maxplus2.all;
LIBRARY ieee;
USE ieee.std_logic_1164.all; 
USE ieee.std_logic_unsigned.all; 

entity Timer is
port (
 opcode: IN std_logic_vector (3 downto 0);
 data: IN std_logic_vector (7 downto 0);
 clock: In std_logic;
 result: OUT std_logic_vector(7 downto 0);
 flag: OUT std_logic);
end Timer;